// Top Package for MNIST Accelerator Core
package core_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    
    
endpackage