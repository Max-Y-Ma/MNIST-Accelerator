`define DATA_WIDTH (32)
`define INTEGER_WIDTH (17)
`define DECIMAL_WIDTH (`DATA_WIDTH - `INTEGER_WIDTH)
`define LAYER1_WIDTH (784)
`define LAYER2_WIDTH (20)
`define LAYER3_WIDTH (20)
`define LAYER4_WIDTH (10)
`define IMG_WIDTH (28)
`define IMG_HEIGHT (28)
`define TEST_DATA_FILE_PATH ("../../../data/mnist_test.csv")
`define TEST_SAMPLES (500)